library verilog;
use verilog.vl_types.all;
entity lab_7_vlg_vec_tst is
end lab_7_vlg_vec_tst;
