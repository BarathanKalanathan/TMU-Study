library verilog;
use verilog.vl_types.all;
entity pc_comb_ckt_ex2_vlg_vec_tst is
end pc_comb_ckt_ex2_vlg_vec_tst;
